`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:23:02 11/13/2020 
// Design Name: 
// Module Name:    half_adder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
//half adder created for 16 bit ripple carry adder
module half_adder(sum, carry, A, B);
  input A,B;
  output sum, carry;
  xor (sum, A, B);
  and (carry, A, B);
endmodule
